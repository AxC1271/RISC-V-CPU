library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- this is the top module of the CPU where all the modules
-- get connected to be fully functional
entity riscv_processor is
  port (

  );

end riscv_processor;

architecture Behavioral of riscv_process is
begin
  
end Behavioral;
