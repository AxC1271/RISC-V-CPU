entity seven_seg_mux is
  port (
  );
end seven_seg_mux;

architecture Behavioral of seven_seg_mux is
begin
end Behavioral;
