library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- seven seg display driver for the basys3 fpga board

entity seven_seg_mux is
  port (
  );
end seven_seg_mux;

architecture Behavioral of seven_seg_mux is
begin
end Behavioral;
