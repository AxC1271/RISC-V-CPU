entity riscv_processor is
  port (

  );

end riscv_processor;

architecture Behavioral of riscv_process is
begin
  
end Behavioral;
